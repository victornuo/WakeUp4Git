----------------------------------------------------------------------
-- Created by Actel SmartDesign Wed Jan 30 12:10:59 2013
-- Testbench Template
-- This is a basic testbench that instantiates your design with basic 
-- clock and reset pins connected.  If your design has special
-- clock/reset or testbench driver requirements then you should 
-- copy this file and modify it. 
----------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;

entity testbench is
end testbench;

architecture behavioral of testbench is

    constant SYSCLK_PERIOD : time := 100 ns;

    signal SYSCLK : std_logic := '0';
    signal NSYSRESET : std_logic := '0';

    component WuPu
        -- ports
        port( 
            -- Inputs
            clk : in std_logic;
            RX : in std_logic;
            RST : in std_logic;
            Flash_Freeze_N : in std_logic;

            -- Outputs
            RESETZB : out std_logic;
            RX_OUT : out std_logic;
            AddOKflag : out std_logic;
            bit_error : out std_logic;
            NewMsg : out std_logic;
            dout : out std_logic;
            new_data : out std_logic;
            d_hk : out std_logic

            -- Inouts

        );
    end component;

begin

    process
        variable vhdl_initial : BOOLEAN := TRUE;

    begin
        if ( vhdl_initial ) then
            -- Assert Reset
            NSYSRESET <= '0';
            wait for ( SYSCLK_PERIOD * 10 );
            
            NSYSRESET <= '1';
            wait;
        end if;
    end process;

    -- 10MHz Clock Driver
    SYSCLK <= not SYSCLK after (SYSCLK_PERIOD / 2.0 );

    -- Instantiate Unit Under Test:  WuPu
    WuPu_0 : WuPu
        -- port map
        port map( 
            -- Inputs
            clk => SYSCLK,
            RX => '0',
            RST => NSYSRESET,
            Flash_Freeze_N => '0',

            -- Outputs
            RESETZB =>  open,
            RX_OUT =>  open,
            AddOKflag =>  open,
            bit_error =>  open,
            NewMsg =>  open,
            dout =>  open,
            new_data =>  open,
            d_hk =>  open

            -- Inouts

        );

end behavioral;

